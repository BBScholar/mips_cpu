

module register_file_logic(
    rs, rt, rd,
    hi, lo, pc_p4, 
    read_data1, read_data2    
);

    register_file rf();

endmodule