

module dff(d, clk, q, qb);

    

endmodule